[HTMLEFS][1][MiniCog][Enterprise, VMC , Test][Mini-Cog; Created by Derry Everson 06/13/2019][MiniCog][//localserver/EncounterForms/HtmlForms/MiniCog/minicog.html][Arial]
