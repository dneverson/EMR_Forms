[HTMLEFS][1][HCCSearch][Enterprise, VMC , Test][HCCSearch; Created by Derry Everson 11/05/2018][HCCSearch][//localserver/EncounterForms/HtmlForms/HCCSearch/index.html][Arial]
