[HTMLEFS][1][In Home Visit][Enterprise, VMC , Test][In Home Encounter; Created by Derry Everson 11/25/2019][In Home Visit][//localserver/EncounterForms/HtmlForms/HomeCareManagement/HomeEncounter.html][Arial]
