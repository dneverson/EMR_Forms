[HTMLEFS][1][QMAF][Enterprise, VMC , Test][QMAF; Created by Robin W. 2016][QMAF][//localserver/EncounterForms/HtmlForms/QualityMeasures/QualityMeasures.html][Arial]
