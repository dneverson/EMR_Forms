[HTMLEFS][1][VBR][Enterprise, VMC , Test][Value Based Revenue; Created by Derry Everson 06/13/2019][VBR][//localserver/EncounterForms/HtmlForms/VBR/vbr.html][Arial]
