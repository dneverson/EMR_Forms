[HTMLEFS][1][Referrals][Enterprise, VMC , Test][Referrals; Created by Robin W. 2017][Referrals][//localserver/EncounterForms/HtmlForms/Referrals/index.html][Arial]
